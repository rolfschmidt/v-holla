module holla

import sqlite

pub fn sqlite_example() bool {
    db := sqlite.connect('holla.db') or {
        panic('driver init failed:$err')
    }

    return true
}