module holla

//fn test_example() {
//    assert postgresql_example() == true
//}