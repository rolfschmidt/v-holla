module holla

//fn test_example() {
//    assert sqlite_example() == true
//}