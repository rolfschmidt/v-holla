module holla

fn test_example() {
    assert mysql_example() == true
}